/////////////////// Please synthesize this RO with lvt library /////////////////// 
/////////////////// This RO contains 383 stages /////////////////// 

`timescale 1ps / 100fs

module RO_inv_slvt(
input wire i_Enable,
input wire i_Sel,
output wire o_RO_out
);

/////////////////// Define wires between inverters ///////////////////
wire [382:0] w_inv_Conn;

NAND3_X2R_A9PP84TSL_C14 U0(
.A(i_Enable),
.B(i_Sel),
.C(o_RO_out),
.Y(w_inv_Conn[0])
);

inv_slvt U1(
.in(w_inv_Conn[0]),
.out(w_inv_Conn[1])
);

inv_slvt U2(
.in(w_inv_Conn[1]),
.out(w_inv_Conn[2])
);

inv_slvt U3(
.in(w_inv_Conn[2]),
.out(w_inv_Conn[3])
);

inv_slvt U4(
.in(w_inv_Conn[3]),
.out(w_inv_Conn[4])
);

inv_slvt U5(
.in(w_inv_Conn[4]),
.out(w_inv_Conn[5])
);

inv_slvt U6(
.in(w_inv_Conn[5]),
.out(w_inv_Conn[6])
);

inv_slvt U7(
.in(w_inv_Conn[6]),
.out(w_inv_Conn[7])
);

inv_slvt U8(
.in(w_inv_Conn[7]),
.out(w_inv_Conn[8])
);

inv_slvt U9(
.in(w_inv_Conn[8]),
.out(w_inv_Conn[9])
);

inv_slvt U10(
.in(w_inv_Conn[9]),
.out(w_inv_Conn[10])
);

inv_slvt U11(
.in(w_inv_Conn[10]),
.out(w_inv_Conn[11])
);

inv_slvt U12(
.in(w_inv_Conn[11]),
.out(w_inv_Conn[12])
);

inv_slvt U13(
.in(w_inv_Conn[12]),
.out(w_inv_Conn[13])
);

inv_slvt U14(
.in(w_inv_Conn[13]),
.out(w_inv_Conn[14])
);

inv_slvt U15(
.in(w_inv_Conn[14]),
.out(w_inv_Conn[15])
);

inv_slvt U16(
.in(w_inv_Conn[15]),
.out(w_inv_Conn[16])
);

inv_slvt U17(
.in(w_inv_Conn[16]),
.out(w_inv_Conn[17])
);

inv_slvt U18(
.in(w_inv_Conn[17]),
.out(w_inv_Conn[18])
);

inv_slvt U19(
.in(w_inv_Conn[18]),
.out(w_inv_Conn[19])
);

inv_slvt U20(
.in(w_inv_Conn[19]),
.out(w_inv_Conn[20])
);

inv_slvt U21(
.in(w_inv_Conn[20]),
.out(w_inv_Conn[21])
);

inv_slvt U22(
.in(w_inv_Conn[21]),
.out(w_inv_Conn[22])
);

inv_slvt U23(
.in(w_inv_Conn[22]),
.out(w_inv_Conn[23])
);

inv_slvt U24(
.in(w_inv_Conn[23]),
.out(w_inv_Conn[24])
);

inv_slvt U25(
.in(w_inv_Conn[24]),
.out(w_inv_Conn[25])
);

inv_slvt U26(
.in(w_inv_Conn[25]),
.out(w_inv_Conn[26])
);

inv_slvt U27(
.in(w_inv_Conn[26]),
.out(w_inv_Conn[27])
);

inv_slvt U28(
.in(w_inv_Conn[27]),
.out(w_inv_Conn[28])
);

inv_slvt U29(
.in(w_inv_Conn[28]),
.out(w_inv_Conn[29])
);

inv_slvt U30(
.in(w_inv_Conn[29]),
.out(w_inv_Conn[30])
);

inv_slvt U31(
.in(w_inv_Conn[30]),
.out(w_inv_Conn[31])
);

inv_slvt U32(
.in(w_inv_Conn[31]),
.out(w_inv_Conn[32])
);

inv_slvt U33(
.in(w_inv_Conn[32]),
.out(w_inv_Conn[33])
);

inv_slvt U34(
.in(w_inv_Conn[33]),
.out(w_inv_Conn[34])
);

inv_slvt U35(
.in(w_inv_Conn[34]),
.out(w_inv_Conn[35])
);

inv_slvt U36(
.in(w_inv_Conn[35]),
.out(w_inv_Conn[36])
);

inv_slvt U37(
.in(w_inv_Conn[36]),
.out(w_inv_Conn[37])
);

inv_slvt U38(
.in(w_inv_Conn[37]),
.out(w_inv_Conn[38])
);

inv_slvt U39(
.in(w_inv_Conn[38]),
.out(w_inv_Conn[39])
);

inv_slvt U40(
.in(w_inv_Conn[39]),
.out(w_inv_Conn[40])
);

inv_slvt U41(
.in(w_inv_Conn[40]),
.out(w_inv_Conn[41])
);

inv_slvt U42(
.in(w_inv_Conn[41]),
.out(w_inv_Conn[42])
);

inv_slvt U43(
.in(w_inv_Conn[42]),
.out(w_inv_Conn[43])
);

inv_slvt U44(
.in(w_inv_Conn[43]),
.out(w_inv_Conn[44])
);

inv_slvt U45(
.in(w_inv_Conn[44]),
.out(w_inv_Conn[45])
);

inv_slvt U46(
.in(w_inv_Conn[45]),
.out(w_inv_Conn[46])
);

inv_slvt U47(
.in(w_inv_Conn[46]),
.out(w_inv_Conn[47])
);

inv_slvt U48(
.in(w_inv_Conn[47]),
.out(w_inv_Conn[48])
);

inv_slvt U49(
.in(w_inv_Conn[48]),
.out(w_inv_Conn[49])
);

inv_slvt U50(
.in(w_inv_Conn[49]),
.out(w_inv_Conn[50])
);

inv_slvt U51(
.in(w_inv_Conn[50]),
.out(w_inv_Conn[51])
);

inv_slvt U52(
.in(w_inv_Conn[51]),
.out(w_inv_Conn[52])
);

inv_slvt U53(
.in(w_inv_Conn[52]),
.out(w_inv_Conn[53])
);

inv_slvt U54(
.in(w_inv_Conn[53]),
.out(w_inv_Conn[54])
);

inv_slvt U55(
.in(w_inv_Conn[54]),
.out(w_inv_Conn[55])
);

inv_slvt U56(
.in(w_inv_Conn[55]),
.out(w_inv_Conn[56])
);

inv_slvt U57(
.in(w_inv_Conn[56]),
.out(w_inv_Conn[57])
);

inv_slvt U58(
.in(w_inv_Conn[57]),
.out(w_inv_Conn[58])
);

inv_slvt U59(
.in(w_inv_Conn[58]),
.out(w_inv_Conn[59])
);

inv_slvt U60(
.in(w_inv_Conn[59]),
.out(w_inv_Conn[60])
);

inv_slvt U61(
.in(w_inv_Conn[60]),
.out(w_inv_Conn[61])
);

inv_slvt U62(
.in(w_inv_Conn[61]),
.out(w_inv_Conn[62])
);

inv_slvt U63(
.in(w_inv_Conn[62]),
.out(w_inv_Conn[63])
);

inv_slvt U64(
.in(w_inv_Conn[63]),
.out(w_inv_Conn[64])
);

inv_slvt U65(
.in(w_inv_Conn[64]),
.out(w_inv_Conn[65])
);

inv_slvt U66(
.in(w_inv_Conn[65]),
.out(w_inv_Conn[66])
);

inv_slvt U67(
.in(w_inv_Conn[66]),
.out(w_inv_Conn[67])
);

inv_slvt U68(
.in(w_inv_Conn[67]),
.out(w_inv_Conn[68])
);

inv_slvt U69(
.in(w_inv_Conn[68]),
.out(w_inv_Conn[69])
);

inv_slvt U70(
.in(w_inv_Conn[69]),
.out(w_inv_Conn[70])
);

inv_slvt U71(
.in(w_inv_Conn[70]),
.out(w_inv_Conn[71])
);

inv_slvt U72(
.in(w_inv_Conn[71]),
.out(w_inv_Conn[72])
);

inv_slvt U73(
.in(w_inv_Conn[72]),
.out(w_inv_Conn[73])
);

inv_slvt U74(
.in(w_inv_Conn[73]),
.out(w_inv_Conn[74])
);

inv_slvt U75(
.in(w_inv_Conn[74]),
.out(w_inv_Conn[75])
);

inv_slvt U76(
.in(w_inv_Conn[75]),
.out(w_inv_Conn[76])
);

inv_slvt U77(
.in(w_inv_Conn[76]),
.out(w_inv_Conn[77])
);

inv_slvt U78(
.in(w_inv_Conn[77]),
.out(w_inv_Conn[78])
);

inv_slvt U79(
.in(w_inv_Conn[78]),
.out(w_inv_Conn[79])
);

inv_slvt U80(
.in(w_inv_Conn[79]),
.out(w_inv_Conn[80])
);

inv_slvt U81(
.in(w_inv_Conn[80]),
.out(w_inv_Conn[81])
);

inv_slvt U82(
.in(w_inv_Conn[81]),
.out(w_inv_Conn[82])
);

inv_slvt U83(
.in(w_inv_Conn[82]),
.out(w_inv_Conn[83])
);

inv_slvt U84(
.in(w_inv_Conn[83]),
.out(w_inv_Conn[84])
);

inv_slvt U85(
.in(w_inv_Conn[84]),
.out(w_inv_Conn[85])
);

inv_slvt U86(
.in(w_inv_Conn[85]),
.out(w_inv_Conn[86])
);

inv_slvt U87(
.in(w_inv_Conn[86]),
.out(w_inv_Conn[87])
);

inv_slvt U88(
.in(w_inv_Conn[87]),
.out(w_inv_Conn[88])
);

inv_slvt U89(
.in(w_inv_Conn[88]),
.out(w_inv_Conn[89])
);

inv_slvt U90(
.in(w_inv_Conn[89]),
.out(w_inv_Conn[90])
);

inv_slvt U91(
.in(w_inv_Conn[90]),
.out(w_inv_Conn[91])
);

inv_slvt U92(
.in(w_inv_Conn[91]),
.out(w_inv_Conn[92])
);

inv_slvt U93(
.in(w_inv_Conn[92]),
.out(w_inv_Conn[93])
);

inv_slvt U94(
.in(w_inv_Conn[93]),
.out(w_inv_Conn[94])
);

inv_slvt U95(
.in(w_inv_Conn[94]),
.out(w_inv_Conn[95])
);

inv_slvt U96(
.in(w_inv_Conn[95]),
.out(w_inv_Conn[96])
);

inv_slvt U97(
.in(w_inv_Conn[96]),
.out(w_inv_Conn[97])
);

inv_slvt U98(
.in(w_inv_Conn[97]),
.out(w_inv_Conn[98])
);

inv_slvt U99(
.in(w_inv_Conn[98]),
.out(w_inv_Conn[99])
);

inv_slvt U100(
.in(w_inv_Conn[99]),
.out(w_inv_Conn[100])
);

inv_slvt U101(
.in(w_inv_Conn[100]),
.out(w_inv_Conn[101])
);

inv_slvt U102(
.in(w_inv_Conn[101]),
.out(w_inv_Conn[102])
);

inv_slvt U103(
.in(w_inv_Conn[102]),
.out(w_inv_Conn[103])
);

inv_slvt U104(
.in(w_inv_Conn[103]),
.out(w_inv_Conn[104])
);

inv_slvt U105(
.in(w_inv_Conn[104]),
.out(w_inv_Conn[105])
);

inv_slvt U106(
.in(w_inv_Conn[105]),
.out(w_inv_Conn[106])
);

inv_slvt U107(
.in(w_inv_Conn[106]),
.out(w_inv_Conn[107])
);

inv_slvt U108(
.in(w_inv_Conn[107]),
.out(w_inv_Conn[108])
);

inv_slvt U109(
.in(w_inv_Conn[108]),
.out(w_inv_Conn[109])
);

inv_slvt U110(
.in(w_inv_Conn[109]),
.out(w_inv_Conn[110])
);

inv_slvt U111(
.in(w_inv_Conn[110]),
.out(w_inv_Conn[111])
);

inv_slvt U112(
.in(w_inv_Conn[111]),
.out(w_inv_Conn[112])
);

inv_slvt U113(
.in(w_inv_Conn[112]),
.out(w_inv_Conn[113])
);

inv_slvt U114(
.in(w_inv_Conn[113]),
.out(w_inv_Conn[114])
);

inv_slvt U115(
.in(w_inv_Conn[114]),
.out(w_inv_Conn[115])
);

inv_slvt U116(
.in(w_inv_Conn[115]),
.out(w_inv_Conn[116])
);

inv_slvt U117(
.in(w_inv_Conn[116]),
.out(w_inv_Conn[117])
);

inv_slvt U118(
.in(w_inv_Conn[117]),
.out(w_inv_Conn[118])
);

inv_slvt U119(
.in(w_inv_Conn[118]),
.out(w_inv_Conn[119])
);

inv_slvt U120(
.in(w_inv_Conn[119]),
.out(w_inv_Conn[120])
);

inv_slvt U121(
.in(w_inv_Conn[120]),
.out(w_inv_Conn[121])
);

inv_slvt U122(
.in(w_inv_Conn[121]),
.out(w_inv_Conn[122])
);

inv_slvt U123(
.in(w_inv_Conn[122]),
.out(w_inv_Conn[123])
);

inv_slvt U124(
.in(w_inv_Conn[123]),
.out(w_inv_Conn[124])
);

inv_slvt U125(
.in(w_inv_Conn[124]),
.out(w_inv_Conn[125])
);

inv_slvt U126(
.in(w_inv_Conn[125]),
.out(w_inv_Conn[126])
);

inv_slvt U127(
.in(w_inv_Conn[126]),
.out(w_inv_Conn[127])
);

inv_slvt U128(
.in(w_inv_Conn[127]),
.out(w_inv_Conn[128])
);

inv_slvt U129(
.in(w_inv_Conn[128]),
.out(w_inv_Conn[129])
);

inv_slvt U130(
.in(w_inv_Conn[129]),
.out(w_inv_Conn[130])
);

inv_slvt U131(
.in(w_inv_Conn[130]),
.out(w_inv_Conn[131])
);

inv_slvt U132(
.in(w_inv_Conn[131]),
.out(w_inv_Conn[132])
);

inv_slvt U133(
.in(w_inv_Conn[132]),
.out(w_inv_Conn[133])
);

inv_slvt U134(
.in(w_inv_Conn[133]),
.out(w_inv_Conn[134])
);

inv_slvt U135(
.in(w_inv_Conn[134]),
.out(w_inv_Conn[135])
);

inv_slvt U136(
.in(w_inv_Conn[135]),
.out(w_inv_Conn[136])
);

inv_slvt U137(
.in(w_inv_Conn[136]),
.out(w_inv_Conn[137])
);

inv_slvt U138(
.in(w_inv_Conn[137]),
.out(w_inv_Conn[138])
);

inv_slvt U139(
.in(w_inv_Conn[138]),
.out(w_inv_Conn[139])
);

inv_slvt U140(
.in(w_inv_Conn[139]),
.out(w_inv_Conn[140])
);

inv_slvt U141(
.in(w_inv_Conn[140]),
.out(w_inv_Conn[141])
);

inv_slvt U142(
.in(w_inv_Conn[141]),
.out(w_inv_Conn[142])
);

inv_slvt U143(
.in(w_inv_Conn[142]),
.out(w_inv_Conn[143])
);

inv_slvt U144(
.in(w_inv_Conn[143]),
.out(w_inv_Conn[144])
);

inv_slvt U145(
.in(w_inv_Conn[144]),
.out(w_inv_Conn[145])
);

inv_slvt U146(
.in(w_inv_Conn[145]),
.out(w_inv_Conn[146])
);

inv_slvt U147(
.in(w_inv_Conn[146]),
.out(w_inv_Conn[147])
);

inv_slvt U148(
.in(w_inv_Conn[147]),
.out(w_inv_Conn[148])
);

inv_slvt U149(
.in(w_inv_Conn[148]),
.out(w_inv_Conn[149])
);

inv_slvt U150(
.in(w_inv_Conn[149]),
.out(w_inv_Conn[150])
);

inv_slvt U151(
.in(w_inv_Conn[150]),
.out(w_inv_Conn[151])
);

inv_slvt U152(
.in(w_inv_Conn[151]),
.out(w_inv_Conn[152])
);

inv_slvt U153(
.in(w_inv_Conn[152]),
.out(w_inv_Conn[153])
);

inv_slvt U154(
.in(w_inv_Conn[153]),
.out(w_inv_Conn[154])
);

inv_slvt U155(
.in(w_inv_Conn[154]),
.out(w_inv_Conn[155])
);

inv_slvt U156(
.in(w_inv_Conn[155]),
.out(w_inv_Conn[156])
);

inv_slvt U157(
.in(w_inv_Conn[156]),
.out(w_inv_Conn[157])
);

inv_slvt U158(
.in(w_inv_Conn[157]),
.out(w_inv_Conn[158])
);

inv_slvt U159(
.in(w_inv_Conn[158]),
.out(w_inv_Conn[159])
);

inv_slvt U160(
.in(w_inv_Conn[159]),
.out(w_inv_Conn[160])
);

inv_slvt U161(
.in(w_inv_Conn[160]),
.out(w_inv_Conn[161])
);

inv_slvt U162(
.in(w_inv_Conn[161]),
.out(w_inv_Conn[162])
);

inv_slvt U163(
.in(w_inv_Conn[162]),
.out(w_inv_Conn[163])
);

inv_slvt U164(
.in(w_inv_Conn[163]),
.out(w_inv_Conn[164])
);

inv_slvt U165(
.in(w_inv_Conn[164]),
.out(w_inv_Conn[165])
);

inv_slvt U166(
.in(w_inv_Conn[165]),
.out(w_inv_Conn[166])
);

inv_slvt U167(
.in(w_inv_Conn[166]),
.out(w_inv_Conn[167])
);

inv_slvt U168(
.in(w_inv_Conn[167]),
.out(w_inv_Conn[168])
);

inv_slvt U169(
.in(w_inv_Conn[168]),
.out(w_inv_Conn[169])
);

inv_slvt U170(
.in(w_inv_Conn[169]),
.out(w_inv_Conn[170])
);

inv_slvt U171(
.in(w_inv_Conn[170]),
.out(w_inv_Conn[171])
);

inv_slvt U172(
.in(w_inv_Conn[171]),
.out(w_inv_Conn[172])
);

inv_slvt U173(
.in(w_inv_Conn[172]),
.out(w_inv_Conn[173])
);

inv_slvt U174(
.in(w_inv_Conn[173]),
.out(w_inv_Conn[174])
);

inv_slvt U175(
.in(w_inv_Conn[174]),
.out(w_inv_Conn[175])
);

inv_slvt U176(
.in(w_inv_Conn[175]),
.out(w_inv_Conn[176])
);

inv_slvt U177(
.in(w_inv_Conn[176]),
.out(w_inv_Conn[177])
);

inv_slvt U178(
.in(w_inv_Conn[177]),
.out(w_inv_Conn[178])
);

inv_slvt U179(
.in(w_inv_Conn[178]),
.out(w_inv_Conn[179])
);

inv_slvt U180(
.in(w_inv_Conn[179]),
.out(w_inv_Conn[180])
);

inv_slvt U181(
.in(w_inv_Conn[180]),
.out(w_inv_Conn[181])
);

inv_slvt U182(
.in(w_inv_Conn[181]),
.out(w_inv_Conn[182])
);

inv_slvt U183(
.in(w_inv_Conn[182]),
.out(w_inv_Conn[183])
);

inv_slvt U184(
.in(w_inv_Conn[183]),
.out(w_inv_Conn[184])
);

inv_slvt U185(
.in(w_inv_Conn[184]),
.out(w_inv_Conn[185])
);

inv_slvt U186(
.in(w_inv_Conn[185]),
.out(w_inv_Conn[186])
);

inv_slvt U187(
.in(w_inv_Conn[186]),
.out(w_inv_Conn[187])
);

inv_slvt U188(
.in(w_inv_Conn[187]),
.out(w_inv_Conn[188])
);

inv_slvt U189(
.in(w_inv_Conn[188]),
.out(w_inv_Conn[189])
);

inv_slvt U190(
.in(w_inv_Conn[189]),
.out(w_inv_Conn[190])
);

inv_slvt U191(
.in(w_inv_Conn[190]),
.out(w_inv_Conn[191])
);

inv_slvt U192(
.in(w_inv_Conn[191]),
.out(w_inv_Conn[192])
);

inv_slvt U193(
.in(w_inv_Conn[192]),
.out(w_inv_Conn[193])
);

inv_slvt U194(
.in(w_inv_Conn[193]),
.out(w_inv_Conn[194])
);

inv_slvt U195(
.in(w_inv_Conn[194]),
.out(w_inv_Conn[195])
);

inv_slvt U196(
.in(w_inv_Conn[195]),
.out(w_inv_Conn[196])
);

inv_slvt U197(
.in(w_inv_Conn[196]),
.out(w_inv_Conn[197])
);

inv_slvt U198(
.in(w_inv_Conn[197]),
.out(w_inv_Conn[198])
);

inv_slvt U199(
.in(w_inv_Conn[198]),
.out(w_inv_Conn[199])
);

inv_slvt U200(
.in(w_inv_Conn[199]),
.out(w_inv_Conn[200])
);

inv_slvt U201(
.in(w_inv_Conn[200]),
.out(w_inv_Conn[201])
);

inv_slvt U202(
.in(w_inv_Conn[201]),
.out(w_inv_Conn[202])
);

inv_slvt U203(
.in(w_inv_Conn[202]),
.out(w_inv_Conn[203])
);

inv_slvt U204(
.in(w_inv_Conn[203]),
.out(w_inv_Conn[204])
);

inv_slvt U205(
.in(w_inv_Conn[204]),
.out(w_inv_Conn[205])
);

inv_slvt U206(
.in(w_inv_Conn[205]),
.out(w_inv_Conn[206])
);

inv_slvt U207(
.in(w_inv_Conn[206]),
.out(w_inv_Conn[207])
);

inv_slvt U208(
.in(w_inv_Conn[207]),
.out(w_inv_Conn[208])
);

inv_slvt U209(
.in(w_inv_Conn[208]),
.out(w_inv_Conn[209])
);

inv_slvt U210(
.in(w_inv_Conn[209]),
.out(w_inv_Conn[210])
);

inv_slvt U211(
.in(w_inv_Conn[210]),
.out(w_inv_Conn[211])
);

inv_slvt U212(
.in(w_inv_Conn[211]),
.out(w_inv_Conn[212])
);

inv_slvt U213(
.in(w_inv_Conn[212]),
.out(w_inv_Conn[213])
);

inv_slvt U214(
.in(w_inv_Conn[213]),
.out(w_inv_Conn[214])
);

inv_slvt U215(
.in(w_inv_Conn[214]),
.out(w_inv_Conn[215])
);

inv_slvt U216(
.in(w_inv_Conn[215]),
.out(w_inv_Conn[216])
);

inv_slvt U217(
.in(w_inv_Conn[216]),
.out(w_inv_Conn[217])
);

inv_slvt U218(
.in(w_inv_Conn[217]),
.out(w_inv_Conn[218])
);

inv_slvt U219(
.in(w_inv_Conn[218]),
.out(w_inv_Conn[219])
);

inv_slvt U220(
.in(w_inv_Conn[219]),
.out(w_inv_Conn[220])
);

inv_slvt U221(
.in(w_inv_Conn[220]),
.out(w_inv_Conn[221])
);

inv_slvt U222(
.in(w_inv_Conn[221]),
.out(w_inv_Conn[222])
);

inv_slvt U223(
.in(w_inv_Conn[222]),
.out(w_inv_Conn[223])
);

inv_slvt U224(
.in(w_inv_Conn[223]),
.out(w_inv_Conn[224])
);

inv_slvt U225(
.in(w_inv_Conn[224]),
.out(w_inv_Conn[225])
);

inv_slvt U226(
.in(w_inv_Conn[225]),
.out(w_inv_Conn[226])
);

inv_slvt U227(
.in(w_inv_Conn[226]),
.out(w_inv_Conn[227])
);

inv_slvt U228(
.in(w_inv_Conn[227]),
.out(w_inv_Conn[228])
);

inv_slvt U229(
.in(w_inv_Conn[228]),
.out(w_inv_Conn[229])
);

inv_slvt U230(
.in(w_inv_Conn[229]),
.out(w_inv_Conn[230])
);

inv_slvt U231(
.in(w_inv_Conn[230]),
.out(w_inv_Conn[231])
);

inv_slvt U232(
.in(w_inv_Conn[231]),
.out(w_inv_Conn[232])
);

inv_slvt U233(
.in(w_inv_Conn[232]),
.out(w_inv_Conn[233])
);

inv_slvt U234(
.in(w_inv_Conn[233]),
.out(w_inv_Conn[234])
);

inv_slvt U235(
.in(w_inv_Conn[234]),
.out(w_inv_Conn[235])
);

inv_slvt U236(
.in(w_inv_Conn[235]),
.out(w_inv_Conn[236])
);

inv_slvt U237(
.in(w_inv_Conn[236]),
.out(w_inv_Conn[237])
);

inv_slvt U238(
.in(w_inv_Conn[237]),
.out(w_inv_Conn[238])
);

inv_slvt U239(
.in(w_inv_Conn[238]),
.out(w_inv_Conn[239])
);

inv_slvt U240(
.in(w_inv_Conn[239]),
.out(w_inv_Conn[240])
);

inv_slvt U241(
.in(w_inv_Conn[240]),
.out(w_inv_Conn[241])
);

inv_slvt U242(
.in(w_inv_Conn[241]),
.out(w_inv_Conn[242])
);

inv_slvt U243(
.in(w_inv_Conn[242]),
.out(w_inv_Conn[243])
);

inv_slvt U244(
.in(w_inv_Conn[243]),
.out(w_inv_Conn[244])
);

inv_slvt U245(
.in(w_inv_Conn[244]),
.out(w_inv_Conn[245])
);

inv_slvt U246(
.in(w_inv_Conn[245]),
.out(w_inv_Conn[246])
);

inv_slvt U247(
.in(w_inv_Conn[246]),
.out(w_inv_Conn[247])
);

inv_slvt U248(
.in(w_inv_Conn[247]),
.out(w_inv_Conn[248])
);

inv_slvt U249(
.in(w_inv_Conn[248]),
.out(w_inv_Conn[249])
);

inv_slvt U250(
.in(w_inv_Conn[249]),
.out(w_inv_Conn[250])
);

inv_slvt U251(
.in(w_inv_Conn[250]),
.out(w_inv_Conn[251])
);

inv_slvt U252(
.in(w_inv_Conn[251]),
.out(w_inv_Conn[252])
);

inv_slvt U253(
.in(w_inv_Conn[252]),
.out(w_inv_Conn[253])
);

inv_slvt U254(
.in(w_inv_Conn[253]),
.out(w_inv_Conn[254])
);

inv_slvt U255(
.in(w_inv_Conn[254]),
.out(w_inv_Conn[255])
);

inv_slvt U256(
.in(w_inv_Conn[255]),
.out(w_inv_Conn[256])
);

inv_slvt U257(
.in(w_inv_Conn[256]),
.out(w_inv_Conn[257])
);

inv_slvt U258(
.in(w_inv_Conn[257]),
.out(w_inv_Conn[258])
);

inv_slvt U259(
.in(w_inv_Conn[258]),
.out(w_inv_Conn[259])
);

inv_slvt U260(
.in(w_inv_Conn[259]),
.out(w_inv_Conn[260])
);

inv_slvt U261(
.in(w_inv_Conn[260]),
.out(w_inv_Conn[261])
);

inv_slvt U262(
.in(w_inv_Conn[261]),
.out(w_inv_Conn[262])
);

inv_slvt U263(
.in(w_inv_Conn[262]),
.out(w_inv_Conn[263])
);

inv_slvt U264(
.in(w_inv_Conn[263]),
.out(w_inv_Conn[264])
);

inv_slvt U265(
.in(w_inv_Conn[264]),
.out(w_inv_Conn[265])
);

inv_slvt U266(
.in(w_inv_Conn[265]),
.out(w_inv_Conn[266])
);

inv_slvt U267(
.in(w_inv_Conn[266]),
.out(w_inv_Conn[267])
);

inv_slvt U268(
.in(w_inv_Conn[267]),
.out(w_inv_Conn[268])
);

inv_slvt U269(
.in(w_inv_Conn[268]),
.out(w_inv_Conn[269])
);

inv_slvt U270(
.in(w_inv_Conn[269]),
.out(w_inv_Conn[270])
);

inv_slvt U271(
.in(w_inv_Conn[270]),
.out(w_inv_Conn[271])
);

inv_slvt U272(
.in(w_inv_Conn[271]),
.out(w_inv_Conn[272])
);

inv_slvt U273(
.in(w_inv_Conn[272]),
.out(w_inv_Conn[273])
);

inv_slvt U274(
.in(w_inv_Conn[273]),
.out(w_inv_Conn[274])
);

inv_slvt U275(
.in(w_inv_Conn[274]),
.out(w_inv_Conn[275])
);

inv_slvt U276(
.in(w_inv_Conn[275]),
.out(w_inv_Conn[276])
);

inv_slvt U277(
.in(w_inv_Conn[276]),
.out(w_inv_Conn[277])
);

inv_slvt U278(
.in(w_inv_Conn[277]),
.out(w_inv_Conn[278])
);

inv_slvt U279(
.in(w_inv_Conn[278]),
.out(w_inv_Conn[279])
);

inv_slvt U280(
.in(w_inv_Conn[279]),
.out(w_inv_Conn[280])
);

inv_slvt U281(
.in(w_inv_Conn[280]),
.out(w_inv_Conn[281])
);

inv_slvt U282(
.in(w_inv_Conn[281]),
.out(w_inv_Conn[282])
);

inv_slvt U283(
.in(w_inv_Conn[282]),
.out(w_inv_Conn[283])
);

inv_slvt U284(
.in(w_inv_Conn[283]),
.out(w_inv_Conn[284])
);

inv_slvt U285(
.in(w_inv_Conn[284]),
.out(w_inv_Conn[285])
);

inv_slvt U286(
.in(w_inv_Conn[285]),
.out(w_inv_Conn[286])
);

inv_slvt U287(
.in(w_inv_Conn[286]),
.out(w_inv_Conn[287])
);

inv_slvt U288(
.in(w_inv_Conn[287]),
.out(w_inv_Conn[288])
);

inv_slvt U289(
.in(w_inv_Conn[288]),
.out(w_inv_Conn[289])
);

inv_slvt U290(
.in(w_inv_Conn[289]),
.out(w_inv_Conn[290])
);

inv_slvt U291(
.in(w_inv_Conn[290]),
.out(w_inv_Conn[291])
);

inv_slvt U292(
.in(w_inv_Conn[291]),
.out(w_inv_Conn[292])
);

inv_slvt U293(
.in(w_inv_Conn[292]),
.out(w_inv_Conn[293])
);

inv_slvt U294(
.in(w_inv_Conn[293]),
.out(w_inv_Conn[294])
);

inv_slvt U295(
.in(w_inv_Conn[294]),
.out(w_inv_Conn[295])
);

inv_slvt U296(
.in(w_inv_Conn[295]),
.out(w_inv_Conn[296])
);

inv_slvt U297(
.in(w_inv_Conn[296]),
.out(w_inv_Conn[297])
);

inv_slvt U298(
.in(w_inv_Conn[297]),
.out(w_inv_Conn[298])
);

inv_slvt U299(
.in(w_inv_Conn[298]),
.out(w_inv_Conn[299])
);

inv_slvt U300(
.in(w_inv_Conn[299]),
.out(w_inv_Conn[300])
);

inv_slvt U301(
.in(w_inv_Conn[300]),
.out(w_inv_Conn[301])
);

inv_slvt U302(
.in(w_inv_Conn[301]),
.out(w_inv_Conn[302])
);

inv_slvt U303(
.in(w_inv_Conn[302]),
.out(w_inv_Conn[303])
);

inv_slvt U304(
.in(w_inv_Conn[303]),
.out(w_inv_Conn[304])
);

inv_slvt U305(
.in(w_inv_Conn[304]),
.out(w_inv_Conn[305])
);

inv_slvt U306(
.in(w_inv_Conn[305]),
.out(w_inv_Conn[306])
);

inv_slvt U307(
.in(w_inv_Conn[306]),
.out(w_inv_Conn[307])
);

inv_slvt U308(
.in(w_inv_Conn[307]),
.out(w_inv_Conn[308])
);

inv_slvt U309(
.in(w_inv_Conn[308]),
.out(w_inv_Conn[309])
);

inv_slvt U310(
.in(w_inv_Conn[309]),
.out(w_inv_Conn[310])
);

inv_slvt U311(
.in(w_inv_Conn[310]),
.out(w_inv_Conn[311])
);

inv_slvt U312(
.in(w_inv_Conn[311]),
.out(w_inv_Conn[312])
);

inv_slvt U313(
.in(w_inv_Conn[312]),
.out(w_inv_Conn[313])
);

inv_slvt U314(
.in(w_inv_Conn[313]),
.out(w_inv_Conn[314])
);

inv_slvt U315(
.in(w_inv_Conn[314]),
.out(w_inv_Conn[315])
);

inv_slvt U316(
.in(w_inv_Conn[315]),
.out(w_inv_Conn[316])
);

inv_slvt U317(
.in(w_inv_Conn[316]),
.out(w_inv_Conn[317])
);

inv_slvt U318(
.in(w_inv_Conn[317]),
.out(w_inv_Conn[318])
);

inv_slvt U319(
.in(w_inv_Conn[318]),
.out(w_inv_Conn[319])
);

inv_slvt U320(
.in(w_inv_Conn[319]),
.out(w_inv_Conn[320])
);

inv_slvt U321(
.in(w_inv_Conn[320]),
.out(w_inv_Conn[321])
);

inv_slvt U322(
.in(w_inv_Conn[321]),
.out(w_inv_Conn[322])
);

inv_slvt U323(
.in(w_inv_Conn[322]),
.out(w_inv_Conn[323])
);

inv_slvt U324(
.in(w_inv_Conn[323]),
.out(w_inv_Conn[324])
);

inv_slvt U325(
.in(w_inv_Conn[324]),
.out(w_inv_Conn[325])
);

inv_slvt U326(
.in(w_inv_Conn[325]),
.out(w_inv_Conn[326])
);

inv_slvt U327(
.in(w_inv_Conn[326]),
.out(w_inv_Conn[327])
);

inv_slvt U328(
.in(w_inv_Conn[327]),
.out(w_inv_Conn[328])
);

inv_slvt U329(
.in(w_inv_Conn[328]),
.out(w_inv_Conn[329])
);

inv_slvt U330(
.in(w_inv_Conn[329]),
.out(w_inv_Conn[330])
);

inv_slvt U331(
.in(w_inv_Conn[330]),
.out(w_inv_Conn[331])
);

inv_slvt U332(
.in(w_inv_Conn[331]),
.out(w_inv_Conn[332])
);

inv_slvt U333(
.in(w_inv_Conn[332]),
.out(w_inv_Conn[333])
);

inv_slvt U334(
.in(w_inv_Conn[333]),
.out(w_inv_Conn[334])
);

inv_slvt U335(
.in(w_inv_Conn[334]),
.out(w_inv_Conn[335])
);

inv_slvt U336(
.in(w_inv_Conn[335]),
.out(w_inv_Conn[336])
);

inv_slvt U337(
.in(w_inv_Conn[336]),
.out(w_inv_Conn[337])
);

inv_slvt U338(
.in(w_inv_Conn[337]),
.out(w_inv_Conn[338])
);

inv_slvt U339(
.in(w_inv_Conn[338]),
.out(w_inv_Conn[339])
);

inv_slvt U340(
.in(w_inv_Conn[339]),
.out(w_inv_Conn[340])
);

inv_slvt U341(
.in(w_inv_Conn[340]),
.out(w_inv_Conn[341])
);

inv_slvt U342(
.in(w_inv_Conn[341]),
.out(w_inv_Conn[342])
);

inv_slvt U343(
.in(w_inv_Conn[342]),
.out(w_inv_Conn[343])
);

inv_slvt U344(
.in(w_inv_Conn[343]),
.out(w_inv_Conn[344])
);

inv_slvt U345(
.in(w_inv_Conn[344]),
.out(w_inv_Conn[345])
);

inv_slvt U346(
.in(w_inv_Conn[345]),
.out(w_inv_Conn[346])
);

inv_slvt U347(
.in(w_inv_Conn[346]),
.out(w_inv_Conn[347])
);

inv_slvt U348(
.in(w_inv_Conn[347]),
.out(w_inv_Conn[348])
);

inv_slvt U349(
.in(w_inv_Conn[348]),
.out(w_inv_Conn[349])
);

inv_slvt U350(
.in(w_inv_Conn[349]),
.out(w_inv_Conn[350])
);

inv_slvt U351(
.in(w_inv_Conn[350]),
.out(w_inv_Conn[351])
);

inv_slvt U352(
.in(w_inv_Conn[351]),
.out(w_inv_Conn[352])
);

inv_slvt U353(
.in(w_inv_Conn[352]),
.out(w_inv_Conn[353])
);

inv_slvt U354(
.in(w_inv_Conn[353]),
.out(w_inv_Conn[354])
);

inv_slvt U355(
.in(w_inv_Conn[354]),
.out(w_inv_Conn[355])
);

inv_slvt U356(
.in(w_inv_Conn[355]),
.out(w_inv_Conn[356])
);

inv_slvt U357(
.in(w_inv_Conn[356]),
.out(w_inv_Conn[357])
);

inv_slvt U358(
.in(w_inv_Conn[357]),
.out(w_inv_Conn[358])
);

inv_slvt U359(
.in(w_inv_Conn[358]),
.out(w_inv_Conn[359])
);

inv_slvt U360(
.in(w_inv_Conn[359]),
.out(w_inv_Conn[360])
);

inv_slvt U361(
.in(w_inv_Conn[360]),
.out(w_inv_Conn[361])
);

inv_slvt U362(
.in(w_inv_Conn[361]),
.out(w_inv_Conn[362])
);

inv_slvt U363(
.in(w_inv_Conn[362]),
.out(w_inv_Conn[363])
);

inv_slvt U364(
.in(w_inv_Conn[363]),
.out(w_inv_Conn[364])
);

inv_slvt U365(
.in(w_inv_Conn[364]),
.out(w_inv_Conn[365])
);

inv_slvt U366(
.in(w_inv_Conn[365]),
.out(w_inv_Conn[366])
);

inv_slvt U367(
.in(w_inv_Conn[366]),
.out(w_inv_Conn[367])
);

inv_slvt U368(
.in(w_inv_Conn[367]),
.out(w_inv_Conn[368])
);

inv_slvt U369(
.in(w_inv_Conn[368]),
.out(w_inv_Conn[369])
);

inv_slvt U370(
.in(w_inv_Conn[369]),
.out(w_inv_Conn[370])
);

inv_slvt U371(
.in(w_inv_Conn[370]),
.out(w_inv_Conn[371])
);

inv_slvt U372(
.in(w_inv_Conn[371]),
.out(w_inv_Conn[372])
);

inv_slvt U373(
.in(w_inv_Conn[372]),
.out(w_inv_Conn[373])
);

inv_slvt U374(
.in(w_inv_Conn[373]),
.out(w_inv_Conn[374])
);

inv_slvt U375(
.in(w_inv_Conn[374]),
.out(w_inv_Conn[375])
);

inv_slvt U376(
.in(w_inv_Conn[375]),
.out(w_inv_Conn[376])
);

inv_slvt U377(
.in(w_inv_Conn[376]),
.out(w_inv_Conn[377])
);

inv_slvt U378(
.in(w_inv_Conn[377]),
.out(w_inv_Conn[378])
);

inv_slvt U379(
.in(w_inv_Conn[378]),
.out(w_inv_Conn[379])
);

inv_slvt U380(
.in(w_inv_Conn[379]),
.out(w_inv_Conn[380])
);

inv_slvt U381(
.in(w_inv_Conn[380]),
.out(w_inv_Conn[381])
);

inv_slvt U382(
.in(w_inv_Conn[381]),
.out(o_RO_out)
);

endmodule

module inv_slvt(
input wire in,
output wire out
); 

INVP_X0P5N_A9PP84TSL_C14 U0(
.A(in),
.Y(out)
);

endmodule 

