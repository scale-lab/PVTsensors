/////////////////// Please synthesize this RO with slvt library /////////////////// 
/////////////////// This RO contains 383 stages /////////////////// 

`timescale 1ps / 100fs

module RO_inv_lvt_65(
input wire i_Enable,
input wire i_Sel,
output wire o_RO_out
);

/////////////////// Define wires between inverters ///////////////////
wire [381:0] w_inv_Conn;

// RTL for NAND3 with imaginary delay numbers
// always@(w_inv_Conn[381] or i_Sel or i_Enable)
assign #110 o_RO_out =  ~(w_inv_Conn[381] & i_Sel & i_Enable);

inv_lvt U1(
.in(o_RO_out),
.out(w_inv_Conn[0])
);

inv_lvt U2(
.in(w_inv_Conn[0]),
.out(w_inv_Conn[1])
);

inv_lvt U3(
.in(w_inv_Conn[1]),
.out(w_inv_Conn[2])
);

inv_lvt U4(
.in(w_inv_Conn[2]),
.out(w_inv_Conn[3])
);

inv_lvt U5(
.in(w_inv_Conn[3]),
.out(w_inv_Conn[4])
);

inv_lvt U6(
.in(w_inv_Conn[4]),
.out(w_inv_Conn[5])
);

inv_lvt U7(
.in(w_inv_Conn[5]),
.out(w_inv_Conn[6])
);

inv_lvt U8(
.in(w_inv_Conn[6]),
.out(w_inv_Conn[7])
);

inv_lvt U9(
.in(w_inv_Conn[7]),
.out(w_inv_Conn[8])
);

inv_lvt U10(
.in(w_inv_Conn[8]),
.out(w_inv_Conn[9])
);

inv_lvt U11(
.in(w_inv_Conn[9]),
.out(w_inv_Conn[10])
);

inv_lvt U12(
.in(w_inv_Conn[10]),
.out(w_inv_Conn[11])
);

inv_lvt U13(
.in(w_inv_Conn[11]),
.out(w_inv_Conn[12])
);

inv_lvt U14(
.in(w_inv_Conn[12]),
.out(w_inv_Conn[13])
);

inv_lvt U15(
.in(w_inv_Conn[13]),
.out(w_inv_Conn[14])
);

inv_lvt U16(
.in(w_inv_Conn[14]),
.out(w_inv_Conn[15])
);

inv_lvt U17(
.in(w_inv_Conn[15]),
.out(w_inv_Conn[16])
);

inv_lvt U18(
.in(w_inv_Conn[16]),
.out(w_inv_Conn[17])
);

inv_lvt U19(
.in(w_inv_Conn[17]),
.out(w_inv_Conn[18])
);

inv_lvt U20(
.in(w_inv_Conn[18]),
.out(w_inv_Conn[19])
);

inv_lvt U21(
.in(w_inv_Conn[19]),
.out(w_inv_Conn[20])
);

inv_lvt U22(
.in(w_inv_Conn[20]),
.out(w_inv_Conn[21])
);

inv_lvt U23(
.in(w_inv_Conn[21]),
.out(w_inv_Conn[22])
);

inv_lvt U24(
.in(w_inv_Conn[22]),
.out(w_inv_Conn[23])
);

inv_lvt U25(
.in(w_inv_Conn[23]),
.out(w_inv_Conn[24])
);

inv_lvt U26(
.in(w_inv_Conn[24]),
.out(w_inv_Conn[25])
);

inv_lvt U27(
.in(w_inv_Conn[25]),
.out(w_inv_Conn[26])
);

inv_lvt U28(
.in(w_inv_Conn[26]),
.out(w_inv_Conn[27])
);

inv_lvt U29(
.in(w_inv_Conn[27]),
.out(w_inv_Conn[28])
);

inv_lvt U30(
.in(w_inv_Conn[28]),
.out(w_inv_Conn[29])
);

inv_lvt U31(
.in(w_inv_Conn[29]),
.out(w_inv_Conn[30])
);

inv_lvt U32(
.in(w_inv_Conn[30]),
.out(w_inv_Conn[31])
);

inv_lvt U33(
.in(w_inv_Conn[31]),
.out(w_inv_Conn[32])
);

inv_lvt U34(
.in(w_inv_Conn[32]),
.out(w_inv_Conn[33])
);

inv_lvt U35(
.in(w_inv_Conn[33]),
.out(w_inv_Conn[34])
);

inv_lvt U36(
.in(w_inv_Conn[34]),
.out(w_inv_Conn[35])
);

inv_lvt U37(
.in(w_inv_Conn[35]),
.out(w_inv_Conn[36])
);

inv_lvt U38(
.in(w_inv_Conn[36]),
.out(w_inv_Conn[37])
);

inv_lvt U39(
.in(w_inv_Conn[37]),
.out(w_inv_Conn[38])
);

inv_lvt U40(
.in(w_inv_Conn[38]),
.out(w_inv_Conn[39])
);

inv_lvt U41(
.in(w_inv_Conn[39]),
.out(w_inv_Conn[40])
);

inv_lvt U42(
.in(w_inv_Conn[40]),
.out(w_inv_Conn[41])
);

inv_lvt U43(
.in(w_inv_Conn[41]),
.out(w_inv_Conn[42])
);

inv_lvt U44(
.in(w_inv_Conn[42]),
.out(w_inv_Conn[43])
);

inv_lvt U45(
.in(w_inv_Conn[43]),
.out(w_inv_Conn[44])
);

inv_lvt U46(
.in(w_inv_Conn[44]),
.out(w_inv_Conn[45])
);

inv_lvt U47(
.in(w_inv_Conn[45]),
.out(w_inv_Conn[46])
);

inv_lvt U48(
.in(w_inv_Conn[46]),
.out(w_inv_Conn[47])
);

inv_lvt U49(
.in(w_inv_Conn[47]),
.out(w_inv_Conn[48])
);

inv_lvt U50(
.in(w_inv_Conn[48]),
.out(w_inv_Conn[49])
);

inv_lvt U51(
.in(w_inv_Conn[49]),
.out(w_inv_Conn[50])
);

inv_lvt U52(
.in(w_inv_Conn[50]),
.out(w_inv_Conn[51])
);

inv_lvt U53(
.in(w_inv_Conn[51]),
.out(w_inv_Conn[52])
);

inv_lvt U54(
.in(w_inv_Conn[52]),
.out(w_inv_Conn[53])
);

inv_lvt U55(
.in(w_inv_Conn[53]),
.out(w_inv_Conn[54])
);

inv_lvt U56(
.in(w_inv_Conn[54]),
.out(w_inv_Conn[55])
);

inv_lvt U57(
.in(w_inv_Conn[55]),
.out(w_inv_Conn[56])
);

inv_lvt U58(
.in(w_inv_Conn[56]),
.out(w_inv_Conn[57])
);

inv_lvt U59(
.in(w_inv_Conn[57]),
.out(w_inv_Conn[58])
);

inv_lvt U60(
.in(w_inv_Conn[58]),
.out(w_inv_Conn[59])
);

inv_lvt U61(
.in(w_inv_Conn[59]),
.out(w_inv_Conn[60])
);

inv_lvt U62(
.in(w_inv_Conn[60]),
.out(w_inv_Conn[61])
);

inv_lvt U63(
.in(w_inv_Conn[61]),
.out(w_inv_Conn[62])
);

inv_lvt U64(
.in(w_inv_Conn[62]),
.out(w_inv_Conn[63])
);

inv_lvt U65(
.in(w_inv_Conn[63]),
.out(w_inv_Conn[64])
);

inv_lvt U66(
.in(w_inv_Conn[64]),
.out(w_inv_Conn[65])
);

inv_lvt U67(
.in(w_inv_Conn[65]),
.out(w_inv_Conn[66])
);

inv_lvt U68(
.in(w_inv_Conn[66]),
.out(w_inv_Conn[67])
);

inv_lvt U69(
.in(w_inv_Conn[67]),
.out(w_inv_Conn[68])
);

inv_lvt U70(
.in(w_inv_Conn[68]),
.out(w_inv_Conn[69])
);

inv_lvt U71(
.in(w_inv_Conn[69]),
.out(w_inv_Conn[70])
);

inv_lvt U72(
.in(w_inv_Conn[70]),
.out(w_inv_Conn[71])
);

inv_lvt U73(
.in(w_inv_Conn[71]),
.out(w_inv_Conn[72])
);

inv_lvt U74(
.in(w_inv_Conn[72]),
.out(w_inv_Conn[73])
);

inv_lvt U75(
.in(w_inv_Conn[73]),
.out(w_inv_Conn[74])
);

inv_lvt U76(
.in(w_inv_Conn[74]),
.out(w_inv_Conn[75])
);

inv_lvt U77(
.in(w_inv_Conn[75]),
.out(w_inv_Conn[76])
);

inv_lvt U78(
.in(w_inv_Conn[76]),
.out(w_inv_Conn[77])
);

inv_lvt U79(
.in(w_inv_Conn[77]),
.out(w_inv_Conn[78])
);

inv_lvt U80(
.in(w_inv_Conn[78]),
.out(w_inv_Conn[79])
);

inv_lvt U81(
.in(w_inv_Conn[79]),
.out(w_inv_Conn[80])
);

inv_lvt U82(
.in(w_inv_Conn[80]),
.out(w_inv_Conn[81])
);

inv_lvt U83(
.in(w_inv_Conn[81]),
.out(w_inv_Conn[82])
);

inv_lvt U84(
.in(w_inv_Conn[82]),
.out(w_inv_Conn[83])
);

inv_lvt U85(
.in(w_inv_Conn[83]),
.out(w_inv_Conn[84])
);

inv_lvt U86(
.in(w_inv_Conn[84]),
.out(w_inv_Conn[85])
);

inv_lvt U87(
.in(w_inv_Conn[85]),
.out(w_inv_Conn[86])
);

inv_lvt U88(
.in(w_inv_Conn[86]),
.out(w_inv_Conn[87])
);

inv_lvt U89(
.in(w_inv_Conn[87]),
.out(w_inv_Conn[88])
);

inv_lvt U90(
.in(w_inv_Conn[88]),
.out(w_inv_Conn[89])
);

inv_lvt U91(
.in(w_inv_Conn[89]),
.out(w_inv_Conn[90])
);

inv_lvt U92(
.in(w_inv_Conn[90]),
.out(w_inv_Conn[91])
);

inv_lvt U93(
.in(w_inv_Conn[91]),
.out(w_inv_Conn[92])
);

inv_lvt U94(
.in(w_inv_Conn[92]),
.out(w_inv_Conn[93])
);

inv_lvt U95(
.in(w_inv_Conn[93]),
.out(w_inv_Conn[94])
);

inv_lvt U96(
.in(w_inv_Conn[94]),
.out(w_inv_Conn[95])
);

inv_lvt U97(
.in(w_inv_Conn[95]),
.out(w_inv_Conn[96])
);

inv_lvt U98(
.in(w_inv_Conn[96]),
.out(w_inv_Conn[97])
);

inv_lvt U99(
.in(w_inv_Conn[97]),
.out(w_inv_Conn[98])
);

inv_lvt U100(
.in(w_inv_Conn[98]),
.out(w_inv_Conn[99])
);

inv_lvt U101(
.in(w_inv_Conn[99]),
.out(w_inv_Conn[100])
);

inv_lvt U102(
.in(w_inv_Conn[100]),
.out(w_inv_Conn[101])
);

inv_lvt U103(
.in(w_inv_Conn[101]),
.out(w_inv_Conn[102])
);

inv_lvt U104(
.in(w_inv_Conn[102]),
.out(w_inv_Conn[103])
);

inv_lvt U105(
.in(w_inv_Conn[103]),
.out(w_inv_Conn[104])
);

inv_lvt U106(
.in(w_inv_Conn[104]),
.out(w_inv_Conn[105])
);

inv_lvt U107(
.in(w_inv_Conn[105]),
.out(w_inv_Conn[106])
);

inv_lvt U108(
.in(w_inv_Conn[106]),
.out(w_inv_Conn[107])
);

inv_lvt U109(
.in(w_inv_Conn[107]),
.out(w_inv_Conn[108])
);

inv_lvt U110(
.in(w_inv_Conn[108]),
.out(w_inv_Conn[109])
);

inv_lvt U111(
.in(w_inv_Conn[109]),
.out(w_inv_Conn[110])
);

inv_lvt U112(
.in(w_inv_Conn[110]),
.out(w_inv_Conn[111])
);

inv_lvt U113(
.in(w_inv_Conn[111]),
.out(w_inv_Conn[112])
);

inv_lvt U114(
.in(w_inv_Conn[112]),
.out(w_inv_Conn[113])
);

inv_lvt U115(
.in(w_inv_Conn[113]),
.out(w_inv_Conn[114])
);

inv_lvt U116(
.in(w_inv_Conn[114]),
.out(w_inv_Conn[115])
);

inv_lvt U117(
.in(w_inv_Conn[115]),
.out(w_inv_Conn[116])
);

inv_lvt U118(
.in(w_inv_Conn[116]),
.out(w_inv_Conn[117])
);

inv_lvt U119(
.in(w_inv_Conn[117]),
.out(w_inv_Conn[118])
);

inv_lvt U120(
.in(w_inv_Conn[118]),
.out(w_inv_Conn[119])
);

inv_lvt U121(
.in(w_inv_Conn[119]),
.out(w_inv_Conn[120])
);

inv_lvt U122(
.in(w_inv_Conn[120]),
.out(w_inv_Conn[121])
);

inv_lvt U123(
.in(w_inv_Conn[121]),
.out(w_inv_Conn[122])
);

inv_lvt U124(
.in(w_inv_Conn[122]),
.out(w_inv_Conn[123])
);

inv_lvt U125(
.in(w_inv_Conn[123]),
.out(w_inv_Conn[124])
);

inv_lvt U126(
.in(w_inv_Conn[124]),
.out(w_inv_Conn[125])
);

inv_lvt U127(
.in(w_inv_Conn[125]),
.out(w_inv_Conn[126])
);

inv_lvt U128(
.in(w_inv_Conn[126]),
.out(w_inv_Conn[127])
);

inv_lvt U129(
.in(w_inv_Conn[127]),
.out(w_inv_Conn[128])
);

inv_lvt U130(
.in(w_inv_Conn[128]),
.out(w_inv_Conn[129])
);

inv_lvt U131(
.in(w_inv_Conn[129]),
.out(w_inv_Conn[130])
);

inv_lvt U132(
.in(w_inv_Conn[130]),
.out(w_inv_Conn[131])
);

inv_lvt U133(
.in(w_inv_Conn[131]),
.out(w_inv_Conn[132])
);

inv_lvt U134(
.in(w_inv_Conn[132]),
.out(w_inv_Conn[133])
);

inv_lvt U135(
.in(w_inv_Conn[133]),
.out(w_inv_Conn[134])
);

inv_lvt U136(
.in(w_inv_Conn[134]),
.out(w_inv_Conn[135])
);

inv_lvt U137(
.in(w_inv_Conn[135]),
.out(w_inv_Conn[136])
);

inv_lvt U138(
.in(w_inv_Conn[136]),
.out(w_inv_Conn[137])
);

inv_lvt U139(
.in(w_inv_Conn[137]),
.out(w_inv_Conn[138])
);

inv_lvt U140(
.in(w_inv_Conn[138]),
.out(w_inv_Conn[139])
);

inv_lvt U141(
.in(w_inv_Conn[139]),
.out(w_inv_Conn[140])
);

inv_lvt U142(
.in(w_inv_Conn[140]),
.out(w_inv_Conn[141])
);

inv_lvt U143(
.in(w_inv_Conn[141]),
.out(w_inv_Conn[142])
);

inv_lvt U144(
.in(w_inv_Conn[142]),
.out(w_inv_Conn[143])
);

inv_lvt U145(
.in(w_inv_Conn[143]),
.out(w_inv_Conn[144])
);

inv_lvt U146(
.in(w_inv_Conn[144]),
.out(w_inv_Conn[145])
);

inv_lvt U147(
.in(w_inv_Conn[145]),
.out(w_inv_Conn[146])
);

inv_lvt U148(
.in(w_inv_Conn[146]),
.out(w_inv_Conn[147])
);

inv_lvt U149(
.in(w_inv_Conn[147]),
.out(w_inv_Conn[148])
);

inv_lvt U150(
.in(w_inv_Conn[148]),
.out(w_inv_Conn[149])
);

inv_lvt U151(
.in(w_inv_Conn[149]),
.out(w_inv_Conn[150])
);

inv_lvt U152(
.in(w_inv_Conn[150]),
.out(w_inv_Conn[151])
);

inv_lvt U153(
.in(w_inv_Conn[151]),
.out(w_inv_Conn[152])
);

inv_lvt U154(
.in(w_inv_Conn[152]),
.out(w_inv_Conn[153])
);

inv_lvt U155(
.in(w_inv_Conn[153]),
.out(w_inv_Conn[154])
);

inv_lvt U156(
.in(w_inv_Conn[154]),
.out(w_inv_Conn[155])
);

inv_lvt U157(
.in(w_inv_Conn[155]),
.out(w_inv_Conn[156])
);

inv_lvt U158(
.in(w_inv_Conn[156]),
.out(w_inv_Conn[157])
);

inv_lvt U159(
.in(w_inv_Conn[157]),
.out(w_inv_Conn[158])
);

inv_lvt U160(
.in(w_inv_Conn[158]),
.out(w_inv_Conn[159])
);

inv_lvt U161(
.in(w_inv_Conn[159]),
.out(w_inv_Conn[160])
);

inv_lvt U162(
.in(w_inv_Conn[160]),
.out(w_inv_Conn[161])
);

inv_lvt U163(
.in(w_inv_Conn[161]),
.out(w_inv_Conn[162])
);

inv_lvt U164(
.in(w_inv_Conn[162]),
.out(w_inv_Conn[163])
);

inv_lvt U165(
.in(w_inv_Conn[163]),
.out(w_inv_Conn[164])
);

inv_lvt U166(
.in(w_inv_Conn[164]),
.out(w_inv_Conn[165])
);

inv_lvt U167(
.in(w_inv_Conn[165]),
.out(w_inv_Conn[166])
);

inv_lvt U168(
.in(w_inv_Conn[166]),
.out(w_inv_Conn[167])
);

inv_lvt U169(
.in(w_inv_Conn[167]),
.out(w_inv_Conn[168])
);

inv_lvt U170(
.in(w_inv_Conn[168]),
.out(w_inv_Conn[169])
);

inv_lvt U171(
.in(w_inv_Conn[169]),
.out(w_inv_Conn[170])
);

inv_lvt U172(
.in(w_inv_Conn[170]),
.out(w_inv_Conn[171])
);

inv_lvt U173(
.in(w_inv_Conn[171]),
.out(w_inv_Conn[172])
);

inv_lvt U174(
.in(w_inv_Conn[172]),
.out(w_inv_Conn[173])
);

inv_lvt U175(
.in(w_inv_Conn[173]),
.out(w_inv_Conn[174])
);

inv_lvt U176(
.in(w_inv_Conn[174]),
.out(w_inv_Conn[175])
);

inv_lvt U177(
.in(w_inv_Conn[175]),
.out(w_inv_Conn[176])
);

inv_lvt U178(
.in(w_inv_Conn[176]),
.out(w_inv_Conn[177])
);

inv_lvt U179(
.in(w_inv_Conn[177]),
.out(w_inv_Conn[178])
);

inv_lvt U180(
.in(w_inv_Conn[178]),
.out(w_inv_Conn[179])
);

inv_lvt U181(
.in(w_inv_Conn[179]),
.out(w_inv_Conn[180])
);

inv_lvt U182(
.in(w_inv_Conn[180]),
.out(w_inv_Conn[181])
);

inv_lvt U183(
.in(w_inv_Conn[181]),
.out(w_inv_Conn[182])
);

inv_lvt U184(
.in(w_inv_Conn[182]),
.out(w_inv_Conn[183])
);

inv_lvt U185(
.in(w_inv_Conn[183]),
.out(w_inv_Conn[184])
);

inv_lvt U186(
.in(w_inv_Conn[184]),
.out(w_inv_Conn[185])
);

inv_lvt U187(
.in(w_inv_Conn[185]),
.out(w_inv_Conn[186])
);

inv_lvt U188(
.in(w_inv_Conn[186]),
.out(w_inv_Conn[187])
);

inv_lvt U189(
.in(w_inv_Conn[187]),
.out(w_inv_Conn[188])
);

inv_lvt U190(
.in(w_inv_Conn[188]),
.out(w_inv_Conn[189])
);

inv_lvt U191(
.in(w_inv_Conn[189]),
.out(w_inv_Conn[190])
);

inv_lvt U192(
.in(w_inv_Conn[190]),
.out(w_inv_Conn[191])
);

inv_lvt U193(
.in(w_inv_Conn[191]),
.out(w_inv_Conn[192])
);

inv_lvt U194(
.in(w_inv_Conn[192]),
.out(w_inv_Conn[193])
);

inv_lvt U195(
.in(w_inv_Conn[193]),
.out(w_inv_Conn[194])
);

inv_lvt U196(
.in(w_inv_Conn[194]),
.out(w_inv_Conn[195])
);

inv_lvt U197(
.in(w_inv_Conn[195]),
.out(w_inv_Conn[196])
);

inv_lvt U198(
.in(w_inv_Conn[196]),
.out(w_inv_Conn[197])
);

inv_lvt U199(
.in(w_inv_Conn[197]),
.out(w_inv_Conn[198])
);

inv_lvt U200(
.in(w_inv_Conn[198]),
.out(w_inv_Conn[199])
);

inv_lvt U201(
.in(w_inv_Conn[199]),
.out(w_inv_Conn[200])
);

inv_lvt U202(
.in(w_inv_Conn[200]),
.out(w_inv_Conn[201])
);

inv_lvt U203(
.in(w_inv_Conn[201]),
.out(w_inv_Conn[202])
);

inv_lvt U204(
.in(w_inv_Conn[202]),
.out(w_inv_Conn[203])
);

inv_lvt U205(
.in(w_inv_Conn[203]),
.out(w_inv_Conn[204])
);

inv_lvt U206(
.in(w_inv_Conn[204]),
.out(w_inv_Conn[205])
);

inv_lvt U207(
.in(w_inv_Conn[205]),
.out(w_inv_Conn[206])
);

inv_lvt U208(
.in(w_inv_Conn[206]),
.out(w_inv_Conn[207])
);

inv_lvt U209(
.in(w_inv_Conn[207]),
.out(w_inv_Conn[208])
);

inv_lvt U210(
.in(w_inv_Conn[208]),
.out(w_inv_Conn[209])
);

inv_lvt U211(
.in(w_inv_Conn[209]),
.out(w_inv_Conn[210])
);

inv_lvt U212(
.in(w_inv_Conn[210]),
.out(w_inv_Conn[211])
);

inv_lvt U213(
.in(w_inv_Conn[211]),
.out(w_inv_Conn[212])
);

inv_lvt U214(
.in(w_inv_Conn[212]),
.out(w_inv_Conn[213])
);

inv_lvt U215(
.in(w_inv_Conn[213]),
.out(w_inv_Conn[214])
);

inv_lvt U216(
.in(w_inv_Conn[214]),
.out(w_inv_Conn[215])
);

inv_lvt U217(
.in(w_inv_Conn[215]),
.out(w_inv_Conn[216])
);

inv_lvt U218(
.in(w_inv_Conn[216]),
.out(w_inv_Conn[217])
);

inv_lvt U219(
.in(w_inv_Conn[217]),
.out(w_inv_Conn[218])
);

inv_lvt U220(
.in(w_inv_Conn[218]),
.out(w_inv_Conn[219])
);

inv_lvt U221(
.in(w_inv_Conn[219]),
.out(w_inv_Conn[220])
);

inv_lvt U222(
.in(w_inv_Conn[220]),
.out(w_inv_Conn[221])
);

inv_lvt U223(
.in(w_inv_Conn[221]),
.out(w_inv_Conn[222])
);

inv_lvt U224(
.in(w_inv_Conn[222]),
.out(w_inv_Conn[223])
);

inv_lvt U225(
.in(w_inv_Conn[223]),
.out(w_inv_Conn[224])
);

inv_lvt U226(
.in(w_inv_Conn[224]),
.out(w_inv_Conn[225])
);

inv_lvt U227(
.in(w_inv_Conn[225]),
.out(w_inv_Conn[226])
);

inv_lvt U228(
.in(w_inv_Conn[226]),
.out(w_inv_Conn[227])
);

inv_lvt U229(
.in(w_inv_Conn[227]),
.out(w_inv_Conn[228])
);

inv_lvt U230(
.in(w_inv_Conn[228]),
.out(w_inv_Conn[229])
);

inv_lvt U231(
.in(w_inv_Conn[229]),
.out(w_inv_Conn[230])
);

inv_lvt U232(
.in(w_inv_Conn[230]),
.out(w_inv_Conn[231])
);

inv_lvt U233(
.in(w_inv_Conn[231]),
.out(w_inv_Conn[232])
);

inv_lvt U234(
.in(w_inv_Conn[232]),
.out(w_inv_Conn[233])
);

inv_lvt U235(
.in(w_inv_Conn[233]),
.out(w_inv_Conn[234])
);

inv_lvt U236(
.in(w_inv_Conn[234]),
.out(w_inv_Conn[235])
);

inv_lvt U237(
.in(w_inv_Conn[235]),
.out(w_inv_Conn[236])
);

inv_lvt U238(
.in(w_inv_Conn[236]),
.out(w_inv_Conn[237])
);

inv_lvt U239(
.in(w_inv_Conn[237]),
.out(w_inv_Conn[238])
);

inv_lvt U240(
.in(w_inv_Conn[238]),
.out(w_inv_Conn[239])
);

inv_lvt U241(
.in(w_inv_Conn[239]),
.out(w_inv_Conn[240])
);

inv_lvt U242(
.in(w_inv_Conn[240]),
.out(w_inv_Conn[241])
);

inv_lvt U243(
.in(w_inv_Conn[241]),
.out(w_inv_Conn[242])
);

inv_lvt U244(
.in(w_inv_Conn[242]),
.out(w_inv_Conn[243])
);

inv_lvt U245(
.in(w_inv_Conn[243]),
.out(w_inv_Conn[244])
);

inv_lvt U246(
.in(w_inv_Conn[244]),
.out(w_inv_Conn[245])
);

inv_lvt U247(
.in(w_inv_Conn[245]),
.out(w_inv_Conn[246])
);

inv_lvt U248(
.in(w_inv_Conn[246]),
.out(w_inv_Conn[247])
);

inv_lvt U249(
.in(w_inv_Conn[247]),
.out(w_inv_Conn[248])
);

inv_lvt U250(
.in(w_inv_Conn[248]),
.out(w_inv_Conn[249])
);

inv_lvt U251(
.in(w_inv_Conn[249]),
.out(w_inv_Conn[250])
);

inv_lvt U252(
.in(w_inv_Conn[250]),
.out(w_inv_Conn[251])
);

inv_lvt U253(
.in(w_inv_Conn[251]),
.out(w_inv_Conn[252])
);

inv_lvt U254(
.in(w_inv_Conn[252]),
.out(w_inv_Conn[253])
);

inv_lvt U255(
.in(w_inv_Conn[253]),
.out(w_inv_Conn[254])
);

inv_lvt U256(
.in(w_inv_Conn[254]),
.out(w_inv_Conn[255])
);

inv_lvt U257(
.in(w_inv_Conn[255]),
.out(w_inv_Conn[256])
);

inv_lvt U258(
.in(w_inv_Conn[256]),
.out(w_inv_Conn[257])
);

inv_lvt U259(
.in(w_inv_Conn[257]),
.out(w_inv_Conn[258])
);

inv_lvt U260(
.in(w_inv_Conn[258]),
.out(w_inv_Conn[259])
);

inv_lvt U261(
.in(w_inv_Conn[259]),
.out(w_inv_Conn[260])
);

inv_lvt U262(
.in(w_inv_Conn[260]),
.out(w_inv_Conn[261])
);

inv_lvt U263(
.in(w_inv_Conn[261]),
.out(w_inv_Conn[262])
);

inv_lvt U264(
.in(w_inv_Conn[262]),
.out(w_inv_Conn[263])
);

inv_lvt U265(
.in(w_inv_Conn[263]),
.out(w_inv_Conn[264])
);

inv_lvt U266(
.in(w_inv_Conn[264]),
.out(w_inv_Conn[265])
);

inv_lvt U267(
.in(w_inv_Conn[265]),
.out(w_inv_Conn[266])
);

inv_lvt U268(
.in(w_inv_Conn[266]),
.out(w_inv_Conn[267])
);

inv_lvt U269(
.in(w_inv_Conn[267]),
.out(w_inv_Conn[268])
);

inv_lvt U270(
.in(w_inv_Conn[268]),
.out(w_inv_Conn[269])
);

inv_lvt U271(
.in(w_inv_Conn[269]),
.out(w_inv_Conn[270])
);

inv_lvt U272(
.in(w_inv_Conn[270]),
.out(w_inv_Conn[271])
);

inv_lvt U273(
.in(w_inv_Conn[271]),
.out(w_inv_Conn[272])
);

inv_lvt U274(
.in(w_inv_Conn[272]),
.out(w_inv_Conn[273])
);

inv_lvt U275(
.in(w_inv_Conn[273]),
.out(w_inv_Conn[274])
);

inv_lvt U276(
.in(w_inv_Conn[274]),
.out(w_inv_Conn[275])
);

inv_lvt U277(
.in(w_inv_Conn[275]),
.out(w_inv_Conn[276])
);

inv_lvt U278(
.in(w_inv_Conn[276]),
.out(w_inv_Conn[277])
);

inv_lvt U279(
.in(w_inv_Conn[277]),
.out(w_inv_Conn[278])
);

inv_lvt U280(
.in(w_inv_Conn[278]),
.out(w_inv_Conn[279])
);

inv_lvt U281(
.in(w_inv_Conn[279]),
.out(w_inv_Conn[280])
);

inv_lvt U282(
.in(w_inv_Conn[280]),
.out(w_inv_Conn[281])
);

inv_lvt U283(
.in(w_inv_Conn[281]),
.out(w_inv_Conn[282])
);

inv_lvt U284(
.in(w_inv_Conn[282]),
.out(w_inv_Conn[283])
);

inv_lvt U285(
.in(w_inv_Conn[283]),
.out(w_inv_Conn[284])
);

inv_lvt U286(
.in(w_inv_Conn[284]),
.out(w_inv_Conn[285])
);

inv_lvt U287(
.in(w_inv_Conn[285]),
.out(w_inv_Conn[286])
);

inv_lvt U288(
.in(w_inv_Conn[286]),
.out(w_inv_Conn[287])
);

inv_lvt U289(
.in(w_inv_Conn[287]),
.out(w_inv_Conn[288])
);

inv_lvt U290(
.in(w_inv_Conn[288]),
.out(w_inv_Conn[289])
);

inv_lvt U291(
.in(w_inv_Conn[289]),
.out(w_inv_Conn[290])
);

inv_lvt U292(
.in(w_inv_Conn[290]),
.out(w_inv_Conn[291])
);

inv_lvt U293(
.in(w_inv_Conn[291]),
.out(w_inv_Conn[292])
);

inv_lvt U294(
.in(w_inv_Conn[292]),
.out(w_inv_Conn[293])
);

inv_lvt U295(
.in(w_inv_Conn[293]),
.out(w_inv_Conn[294])
);

inv_lvt U296(
.in(w_inv_Conn[294]),
.out(w_inv_Conn[295])
);

inv_lvt U297(
.in(w_inv_Conn[295]),
.out(w_inv_Conn[296])
);

inv_lvt U298(
.in(w_inv_Conn[296]),
.out(w_inv_Conn[297])
);

inv_lvt U299(
.in(w_inv_Conn[297]),
.out(w_inv_Conn[298])
);

inv_lvt U300(
.in(w_inv_Conn[298]),
.out(w_inv_Conn[299])
);

inv_lvt U301(
.in(w_inv_Conn[299]),
.out(w_inv_Conn[300])
);

inv_lvt U302(
.in(w_inv_Conn[300]),
.out(w_inv_Conn[301])
);

inv_lvt U303(
.in(w_inv_Conn[301]),
.out(w_inv_Conn[302])
);

inv_lvt U304(
.in(w_inv_Conn[302]),
.out(w_inv_Conn[303])
);

inv_lvt U305(
.in(w_inv_Conn[303]),
.out(w_inv_Conn[304])
);

inv_lvt U306(
.in(w_inv_Conn[304]),
.out(w_inv_Conn[305])
);

inv_lvt U307(
.in(w_inv_Conn[305]),
.out(w_inv_Conn[306])
);

inv_lvt U308(
.in(w_inv_Conn[306]),
.out(w_inv_Conn[307])
);

inv_lvt U309(
.in(w_inv_Conn[307]),
.out(w_inv_Conn[308])
);

inv_lvt U310(
.in(w_inv_Conn[308]),
.out(w_inv_Conn[309])
);

inv_lvt U311(
.in(w_inv_Conn[309]),
.out(w_inv_Conn[310])
);

inv_lvt U312(
.in(w_inv_Conn[310]),
.out(w_inv_Conn[311])
);

inv_lvt U313(
.in(w_inv_Conn[311]),
.out(w_inv_Conn[312])
);

inv_lvt U314(
.in(w_inv_Conn[312]),
.out(w_inv_Conn[313])
);

inv_lvt U315(
.in(w_inv_Conn[313]),
.out(w_inv_Conn[314])
);

inv_lvt U316(
.in(w_inv_Conn[314]),
.out(w_inv_Conn[315])
);

inv_lvt U317(
.in(w_inv_Conn[315]),
.out(w_inv_Conn[316])
);

inv_lvt U318(
.in(w_inv_Conn[316]),
.out(w_inv_Conn[317])
);

inv_lvt U319(
.in(w_inv_Conn[317]),
.out(w_inv_Conn[318])
);

inv_lvt U320(
.in(w_inv_Conn[318]),
.out(w_inv_Conn[319])
);

inv_lvt U321(
.in(w_inv_Conn[319]),
.out(w_inv_Conn[320])
);

inv_lvt U322(
.in(w_inv_Conn[320]),
.out(w_inv_Conn[321])
);

inv_lvt U323(
.in(w_inv_Conn[321]),
.out(w_inv_Conn[322])
);

inv_lvt U324(
.in(w_inv_Conn[322]),
.out(w_inv_Conn[323])
);

inv_lvt U325(
.in(w_inv_Conn[323]),
.out(w_inv_Conn[324])
);

inv_lvt U326(
.in(w_inv_Conn[324]),
.out(w_inv_Conn[325])
);

inv_lvt U327(
.in(w_inv_Conn[325]),
.out(w_inv_Conn[326])
);

inv_lvt U328(
.in(w_inv_Conn[326]),
.out(w_inv_Conn[327])
);

inv_lvt U329(
.in(w_inv_Conn[327]),
.out(w_inv_Conn[328])
);

inv_lvt U330(
.in(w_inv_Conn[328]),
.out(w_inv_Conn[329])
);

inv_lvt U331(
.in(w_inv_Conn[329]),
.out(w_inv_Conn[330])
);

inv_lvt U332(
.in(w_inv_Conn[330]),
.out(w_inv_Conn[331])
);

inv_lvt U333(
.in(w_inv_Conn[331]),
.out(w_inv_Conn[332])
);

inv_lvt U334(
.in(w_inv_Conn[332]),
.out(w_inv_Conn[333])
);

inv_lvt U335(
.in(w_inv_Conn[333]),
.out(w_inv_Conn[334])
);

inv_lvt U336(
.in(w_inv_Conn[334]),
.out(w_inv_Conn[335])
);

inv_lvt U337(
.in(w_inv_Conn[335]),
.out(w_inv_Conn[336])
);

inv_lvt U338(
.in(w_inv_Conn[336]),
.out(w_inv_Conn[337])
);

inv_lvt U339(
.in(w_inv_Conn[337]),
.out(w_inv_Conn[338])
);

inv_lvt U340(
.in(w_inv_Conn[338]),
.out(w_inv_Conn[339])
);

inv_lvt U341(
.in(w_inv_Conn[339]),
.out(w_inv_Conn[340])
);

inv_lvt U342(
.in(w_inv_Conn[340]),
.out(w_inv_Conn[341])
);

inv_lvt U343(
.in(w_inv_Conn[341]),
.out(w_inv_Conn[342])
);

inv_lvt U344(
.in(w_inv_Conn[342]),
.out(w_inv_Conn[343])
);

inv_lvt U345(
.in(w_inv_Conn[343]),
.out(w_inv_Conn[344])
);

inv_lvt U346(
.in(w_inv_Conn[344]),
.out(w_inv_Conn[345])
);

inv_lvt U347(
.in(w_inv_Conn[345]),
.out(w_inv_Conn[346])
);

inv_lvt U348(
.in(w_inv_Conn[346]),
.out(w_inv_Conn[347])
);

inv_lvt U349(
.in(w_inv_Conn[347]),
.out(w_inv_Conn[348])
);

inv_lvt U350(
.in(w_inv_Conn[348]),
.out(w_inv_Conn[349])
);

inv_lvt U351(
.in(w_inv_Conn[349]),
.out(w_inv_Conn[350])
);

inv_lvt U352(
.in(w_inv_Conn[350]),
.out(w_inv_Conn[351])
);

inv_lvt U353(
.in(w_inv_Conn[351]),
.out(w_inv_Conn[352])
);

inv_lvt U354(
.in(w_inv_Conn[352]),
.out(w_inv_Conn[353])
);

inv_lvt U355(
.in(w_inv_Conn[353]),
.out(w_inv_Conn[354])
);

inv_lvt U356(
.in(w_inv_Conn[354]),
.out(w_inv_Conn[355])
);

inv_lvt U357(
.in(w_inv_Conn[355]),
.out(w_inv_Conn[356])
);

inv_lvt U358(
.in(w_inv_Conn[356]),
.out(w_inv_Conn[357])
);

inv_lvt U359(
.in(w_inv_Conn[357]),
.out(w_inv_Conn[358])
);

inv_lvt U360(
.in(w_inv_Conn[358]),
.out(w_inv_Conn[359])
);

inv_lvt U361(
.in(w_inv_Conn[359]),
.out(w_inv_Conn[360])
);

inv_lvt U362(
.in(w_inv_Conn[360]),
.out(w_inv_Conn[361])
);

inv_lvt U363(
.in(w_inv_Conn[361]),
.out(w_inv_Conn[362])
);

inv_lvt U364(
.in(w_inv_Conn[362]),
.out(w_inv_Conn[363])
);

inv_lvt U365(
.in(w_inv_Conn[363]),
.out(w_inv_Conn[364])
);

inv_lvt U366(
.in(w_inv_Conn[364]),
.out(w_inv_Conn[365])
);

inv_lvt U367(
.in(w_inv_Conn[365]),
.out(w_inv_Conn[366])
);

inv_lvt U368(
.in(w_inv_Conn[366]),
.out(w_inv_Conn[367])
);

inv_lvt U369(
.in(w_inv_Conn[367]),
.out(w_inv_Conn[368])
);

inv_lvt U370(
.in(w_inv_Conn[368]),
.out(w_inv_Conn[369])
);

inv_lvt U371(
.in(w_inv_Conn[369]),
.out(w_inv_Conn[370])
);

inv_lvt U372(
.in(w_inv_Conn[370]),
.out(w_inv_Conn[371])
);

inv_lvt U373(
.in(w_inv_Conn[371]),
.out(w_inv_Conn[372])
);

inv_lvt U374(
.in(w_inv_Conn[372]),
.out(w_inv_Conn[373])
);

inv_lvt U375(
.in(w_inv_Conn[373]),
.out(w_inv_Conn[374])
);

inv_lvt U376(
.in(w_inv_Conn[374]),
.out(w_inv_Conn[375])
);

inv_lvt U377(
.in(w_inv_Conn[375]),
.out(w_inv_Conn[376])
);

inv_lvt U378(
.in(w_inv_Conn[376]),
.out(w_inv_Conn[377])
);

inv_lvt U379(
.in(w_inv_Conn[377]),
.out(w_inv_Conn[378])
);

inv_lvt U380(
.in(w_inv_Conn[378]),
.out(w_inv_Conn[379])
);

inv_lvt U381(
.in(w_inv_Conn[379]),
.out(w_inv_Conn[380])
);

inv_lvt U382(
.in(w_inv_Conn[380]),
.out(w_inv_Conn[381])
);

endmodule

module inv_lvt(
input wire in,
output wire out
); 

assign #60 out = ~in;

endmodule 

