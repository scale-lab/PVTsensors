VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
  LAYER LEF58_TYPE STRING ;
  LAYER LEF58_ENCLOSURE STRING ;
  LAYER LEF58_SPACINGTABLE STRING ;
  LAYER LEF58_MINIMUMCUT STRING ;
  LAYER LEF58_SPACING STRING ;
  LAYER LEF58_VOLTAGESPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
  LAYER LEF58_WIDTHTABLE STRING ;
  LAYER LEF58_AREA STRING ;
  LAYER LEF58_EOLEXTENSIONSPACING STRING ;
  LAYER LEF58_CUTCLASS STRING ;
  LAYER LEF58_EOLENCLOSURE STRING ;
  LAYER LEF58_MINSTEP STRING ;
  LAYER LEF58_MINWIDTH STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;
LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

MACRO Brown_PVTSensor
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN Brown_PVTSensor 0 0 ;
  SIZE 100 BY 50 ;
  SYMMETRY X Y ;
  SITE sc9mcpp84_14lpp;

  PIN o_SPI_MISO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.788 1.087 102.82 1.119 ;
    END
  END o_SPI_MISO
  PIN i_SPI_MOSI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER K1 ;
        RECT 102.756 50.328 102.82 50.392 ;
    END
  END i_SPI_MOSI
  PIN i_SPI_Clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER K1 ;
        RECT 102.756 31.429 102.82 31.493 ;
    END
  END i_SPI_Clk
  PIN i_SPI_CS_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER K1 ;
        RECT 102.756 30.368 102.82 30.432 ;
    END
  END i_SPI_CS_n
  PIN i_Rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER K1 ;
        RECT 102.756 1.834 102.82 1.898 ;
    END
  END i_Rst_n
  PIN i_CntWin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 67.234 0.586 67.266 0.618 ;
    END
  END i_CntWin
  PIN i_Clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 66.251 0.586 66.283 0.618 ;
    END
  END i_Clk
  PIN A_BGR_PS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER K1 ;
        RECT 2.82 25.414 2.884 25.478 ;
    END
  END A_BGR_PS
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER K1 ;
        RECT 73.349 0.586 73.413 0.65 ;
    END
  END GND
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER K1 ;
        RECT 75.015 0.586 75.079 0.65 ;
    END
  END DVDD
  PIN AVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER K1 ;
        RECT 71.538 50.522 71.602 50.586 ;
    END
  END AVDD
  PROPERTY CatenaDesignType "deviceLevel" ;
END Brown_PVTSensor

END LIBRARY
