/////////// This is the testbench for the Digital VT sensor ///////////
/////////// This is a temperory file, please maek sure to change name ///////////
`timescale 1ps / 100fs 
module Digital_VT_tb_RTL; 

//////////// Delcaring wires & registers ////////////
reg SPI_CLK_En, SPI_CLK_Continuous;
reg RSTLOW_offchip;
reg SPI_MOSI_offchip;
reg SPI_CS_offchip;
reg SPI_CTRL_offchip;
reg ENABLE_DUMMY_RO_offchip;

wire SPI_MISO_PAD;
wire SPI_CLK_PAD;
wire RSTLOW_PAD;
wire SPI_MOSI_PAD;
wire SPI_CS_PAD;
wire SPI_CTRL_PAD;
wire ENABLE_DUMMY_RO_PAD;

assign SPI_CLK_PAD = SPI_CLK_Continuous & SPI_CLK_En;
assign SPI_MOSI_PAD = SPI_MOSI_offchip;
assign RSTLOW_PAD = RSTLOW_offchip;
assign SPI_CS_PAD = SPI_CS_offchip;
assign SPI_CTRL_PAD = SPI_CTRL_offchip;
assign ENABLE_DUMMY_RO_PAD = ENABLE_DUMMY_RO_offchip;

// XXX_PAD for offchip connection
// XXX_UC for microcontroller connection
// SPI_CTRL = 1'b0, the mux chooses the offchip connection, SPI talks through ports of "XXX_PAD"
// SPI_CTRL = 1'b1, the mux chooses the microcontroller connection, SPI talks through ports of "XXX_UC"

//////////// Call TDU top level ////////////
DigitalVTSensor_chip_quadsensors_V8 TDU(
.RSTLOW_PAD(RSTLOW_PAD), 
.SPI_MOSI_PAD(SPI_MOSI_PAD), 
.SPI_CLK_PAD(SPI_CLK_PAD), 
.SPI_CS_PAD(SPI_CS_PAD), 
.ENABLE_DUMMY_RO_PAD(ENABLE_DUMMY_RO_PAD), 
.SPI_CTRL_PAD(SPI_CTRL_PAD), 
.SPI_MISO_PAD(SPI_MISO_PAD), 
.SPI_MOSI_UC(1'b1), 
.SPI_MISO_UC(), 
.SPI_CS_UC(1'b1), 
.SPI_CLK_UC(1'b1) 
);

//////////// testbench ////////////
initial 
begin
    RSTLOW_offchip = 1'b0;
    SPI_CS_offchip = 1'b1;
    SPI_MOSI_offchip = 1'b0;
    SPI_CLK_En = 1'b0;
    SPI_CLK_Continuous = 1'b1;
    ENABLE_DUMMY_RO_offchip = 1'b0;
    SPI_CTRL_offchip = 1'b0;
    #50000 RSTLOW_offchip = 1'b1;      // after 5ns, rst goes low (50n)
    #100000 SPI_CS_offchip = 1'b0;
    #20000 SPI_CLK_En = 1'b1;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #0 SPI_CLK_En = 1'b0;
    #30000 SPI_CLK_En = 1'b0;
    #50000 SPI_CS_offchip = 1'b1;
    #1000000 SPI_CS_offchip = 1'b1;
    #100000 SPI_CS_offchip = 1'b0;
    #20000 SPI_CLK_En = 1'b1;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #0 SPI_CLK_En = 1'b0;
    #30000 SPI_CLK_En = 1'b0;
    #50000 SPI_CS_offchip = 1'b1;
    #1000000 SPI_CS_offchip = 1'b1;
    #0 ENABLE_DUMMY_RO_offchip = 1'b1;
    #0 SPI_CTRL_offchip = 1'b1;
    #100000 SPI_CS_offchip = 1'b0;
    #20000 SPI_CLK_En = 1'b1;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b0;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #20000 SPI_MOSI_offchip = 1'b1;
    #80000 SPI_MOSI_offchip = 1'b0;
    #0 SPI_CLK_En = 1'b0;
    #30000 SPI_CLK_En = 1'b0;
    #50000 SPI_CS_offchip = 1'b1;
    #1000000 SPI_CS_offchip = 1'b1;
end

//////////// clock source ////////////
always 
begin
    #50000 SPI_CLK_Continuous = ~SPI_CLK_Continuous;
end
endmodule
