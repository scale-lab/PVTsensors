`timescale 1ps / 100fs

module Dummy_RO_Top(
input wire i_Enable,
input wire [31:0] i_Sel
);

//////////////// Dummy ROs ////////////////

Dummy_RO_cell D0(
.i_Enable(i_Enable),
.i_Sel(i_Sel[0])
);

Dummy_RO_cell D1(
.i_Enable(i_Enable),
.i_Sel(i_Sel[0])
);

Dummy_RO_cell D2(
.i_Enable(i_Enable),
.i_Sel(i_Sel[0])
);

Dummy_RO_cell D3(
.i_Enable(i_Enable),
.i_Sel(i_Sel[0])
);

Dummy_RO_cell D4(
.i_Enable(i_Enable),
.i_Sel(i_Sel[1])
);

Dummy_RO_cell D5(
.i_Enable(i_Enable),
.i_Sel(i_Sel[1])
);

Dummy_RO_cell D6(
.i_Enable(i_Enable),
.i_Sel(i_Sel[1])
);

Dummy_RO_cell D7(
.i_Enable(i_Enable),
.i_Sel(i_Sel[1])
);

Dummy_RO_cell D8(
.i_Enable(i_Enable),
.i_Sel(i_Sel[2])
);

Dummy_RO_cell D9(
.i_Enable(i_Enable),
.i_Sel(i_Sel[2])
);

Dummy_RO_cell D10(
.i_Enable(i_Enable),
.i_Sel(i_Sel[2])
);

Dummy_RO_cell D11(
.i_Enable(i_Enable),
.i_Sel(i_Sel[2])
);

Dummy_RO_cell D12(
.i_Enable(i_Enable),
.i_Sel(i_Sel[3])
);

Dummy_RO_cell D13(
.i_Enable(i_Enable),
.i_Sel(i_Sel[3])
);

Dummy_RO_cell D14(
.i_Enable(i_Enable),
.i_Sel(i_Sel[3])
);

Dummy_RO_cell D15(
.i_Enable(i_Enable),
.i_Sel(i_Sel[3])
);

Dummy_RO_cell D16(
.i_Enable(i_Enable),
.i_Sel(i_Sel[4])
);

Dummy_RO_cell D17(
.i_Enable(i_Enable),
.i_Sel(i_Sel[4])
);

Dummy_RO_cell D18(
.i_Enable(i_Enable),
.i_Sel(i_Sel[4])
);

Dummy_RO_cell D19(
.i_Enable(i_Enable),
.i_Sel(i_Sel[4])
);

Dummy_RO_cell D20(
.i_Enable(i_Enable),
.i_Sel(i_Sel[5])
);

Dummy_RO_cell D21(
.i_Enable(i_Enable),
.i_Sel(i_Sel[5])
);

Dummy_RO_cell D22(
.i_Enable(i_Enable),
.i_Sel(i_Sel[5])
);

Dummy_RO_cell D23(
.i_Enable(i_Enable),
.i_Sel(i_Sel[5])
);

Dummy_RO_cell D24(
.i_Enable(i_Enable),
.i_Sel(i_Sel[6])
);

Dummy_RO_cell D25(
.i_Enable(i_Enable),
.i_Sel(i_Sel[6])
);

Dummy_RO_cell D26(
.i_Enable(i_Enable),
.i_Sel(i_Sel[6])
);

Dummy_RO_cell D27(
.i_Enable(i_Enable),
.i_Sel(i_Sel[6])
);

Dummy_RO_cell D28(
.i_Enable(i_Enable),
.i_Sel(i_Sel[7])
);

Dummy_RO_cell D29(
.i_Enable(i_Enable),
.i_Sel(i_Sel[7])
);

Dummy_RO_cell D30(
.i_Enable(i_Enable),
.i_Sel(i_Sel[7])
);

Dummy_RO_cell D31(
.i_Enable(i_Enable),
.i_Sel(i_Sel[7])
);

Dummy_RO_cell D32(
.i_Enable(i_Enable),
.i_Sel(i_Sel[8])
);

Dummy_RO_cell D33(
.i_Enable(i_Enable),
.i_Sel(i_Sel[8])
);

Dummy_RO_cell D34(
.i_Enable(i_Enable),
.i_Sel(i_Sel[8])
);

Dummy_RO_cell D35(
.i_Enable(i_Enable),
.i_Sel(i_Sel[8])
);

Dummy_RO_cell D36(
.i_Enable(i_Enable),
.i_Sel(i_Sel[9])
);

Dummy_RO_cell D37(
.i_Enable(i_Enable),
.i_Sel(i_Sel[9])
);

Dummy_RO_cell D38(
.i_Enable(i_Enable),
.i_Sel(i_Sel[9])
);

Dummy_RO_cell D39(
.i_Enable(i_Enable),
.i_Sel(i_Sel[9])
);

Dummy_RO_cell D40(
.i_Enable(i_Enable),
.i_Sel(i_Sel[10])
);

Dummy_RO_cell D41(
.i_Enable(i_Enable),
.i_Sel(i_Sel[10])
);

Dummy_RO_cell D42(
.i_Enable(i_Enable),
.i_Sel(i_Sel[10])
);

Dummy_RO_cell D43(
.i_Enable(i_Enable),
.i_Sel(i_Sel[10])
);

Dummy_RO_cell D44(
.i_Enable(i_Enable),
.i_Sel(i_Sel[11])
);

Dummy_RO_cell D45(
.i_Enable(i_Enable),
.i_Sel(i_Sel[11])
);

Dummy_RO_cell D46(
.i_Enable(i_Enable),
.i_Sel(i_Sel[11])
);

Dummy_RO_cell D47(
.i_Enable(i_Enable),
.i_Sel(i_Sel[11])
);

Dummy_RO_cell D48(
.i_Enable(i_Enable),
.i_Sel(i_Sel[12])
);

Dummy_RO_cell D49(
.i_Enable(i_Enable),
.i_Sel(i_Sel[12])
);

Dummy_RO_cell D50(
.i_Enable(i_Enable),
.i_Sel(i_Sel[12])
);

Dummy_RO_cell D51(
.i_Enable(i_Enable),
.i_Sel(i_Sel[12])
);

Dummy_RO_cell D52(
.i_Enable(i_Enable),
.i_Sel(i_Sel[13])
);

Dummy_RO_cell D53(
.i_Enable(i_Enable),
.i_Sel(i_Sel[13])
);

Dummy_RO_cell D54(
.i_Enable(i_Enable),
.i_Sel(i_Sel[13])
);

Dummy_RO_cell D55(
.i_Enable(i_Enable),
.i_Sel(i_Sel[13])
);

Dummy_RO_cell D56(
.i_Enable(i_Enable),
.i_Sel(i_Sel[14])
);

Dummy_RO_cell D57(
.i_Enable(i_Enable),
.i_Sel(i_Sel[14])
);

Dummy_RO_cell D58(
.i_Enable(i_Enable),
.i_Sel(i_Sel[14])
);

Dummy_RO_cell D59(
.i_Enable(i_Enable),
.i_Sel(i_Sel[14])
);

Dummy_RO_cell D60(
.i_Enable(i_Enable),
.i_Sel(i_Sel[15])
);

Dummy_RO_cell D61(
.i_Enable(i_Enable),
.i_Sel(i_Sel[15])
);

Dummy_RO_cell D62(
.i_Enable(i_Enable),
.i_Sel(i_Sel[15])
);

Dummy_RO_cell D63(
.i_Enable(i_Enable),
.i_Sel(i_Sel[15])
);

Dummy_RO_cell D64(
.i_Enable(i_Enable),
.i_Sel(i_Sel[16])
);

Dummy_RO_cell D65(
.i_Enable(i_Enable),
.i_Sel(i_Sel[16])
);

Dummy_RO_cell D66(
.i_Enable(i_Enable),
.i_Sel(i_Sel[16])
);

Dummy_RO_cell D67(
.i_Enable(i_Enable),
.i_Sel(i_Sel[16])
);

Dummy_RO_cell D68(
.i_Enable(i_Enable),
.i_Sel(i_Sel[17])
);

Dummy_RO_cell D69(
.i_Enable(i_Enable),
.i_Sel(i_Sel[17])
);

Dummy_RO_cell D70(
.i_Enable(i_Enable),
.i_Sel(i_Sel[17])
);

Dummy_RO_cell D71(
.i_Enable(i_Enable),
.i_Sel(i_Sel[17])
);

Dummy_RO_cell D72(
.i_Enable(i_Enable),
.i_Sel(i_Sel[18])
);

Dummy_RO_cell D73(
.i_Enable(i_Enable),
.i_Sel(i_Sel[18])
);

Dummy_RO_cell D74(
.i_Enable(i_Enable),
.i_Sel(i_Sel[18])
);

Dummy_RO_cell D75(
.i_Enable(i_Enable),
.i_Sel(i_Sel[18])
);

Dummy_RO_cell D76(
.i_Enable(i_Enable),
.i_Sel(i_Sel[19])
);

Dummy_RO_cell D77(
.i_Enable(i_Enable),
.i_Sel(i_Sel[19])
);

Dummy_RO_cell D78(
.i_Enable(i_Enable),
.i_Sel(i_Sel[19])
);

Dummy_RO_cell D79(
.i_Enable(i_Enable),
.i_Sel(i_Sel[19])
);

Dummy_RO_cell D80(
.i_Enable(i_Enable),
.i_Sel(i_Sel[20])
);

Dummy_RO_cell D81(
.i_Enable(i_Enable),
.i_Sel(i_Sel[20])
);

Dummy_RO_cell D82(
.i_Enable(i_Enable),
.i_Sel(i_Sel[20])
);

Dummy_RO_cell D83(
.i_Enable(i_Enable),
.i_Sel(i_Sel[20])
);

Dummy_RO_cell D84(
.i_Enable(i_Enable),
.i_Sel(i_Sel[21])
);

Dummy_RO_cell D85(
.i_Enable(i_Enable),
.i_Sel(i_Sel[21])
);

Dummy_RO_cell D86(
.i_Enable(i_Enable),
.i_Sel(i_Sel[21])
);

Dummy_RO_cell D87(
.i_Enable(i_Enable),
.i_Sel(i_Sel[21])
);

Dummy_RO_cell D88(
.i_Enable(i_Enable),
.i_Sel(i_Sel[22])
);

Dummy_RO_cell D89(
.i_Enable(i_Enable),
.i_Sel(i_Sel[22])
);

Dummy_RO_cell D90(
.i_Enable(i_Enable),
.i_Sel(i_Sel[22])
);

Dummy_RO_cell D91(
.i_Enable(i_Enable),
.i_Sel(i_Sel[22])
);

Dummy_RO_cell D92(
.i_Enable(i_Enable),
.i_Sel(i_Sel[23])
);

Dummy_RO_cell D93(
.i_Enable(i_Enable),
.i_Sel(i_Sel[23])
);

Dummy_RO_cell D94(
.i_Enable(i_Enable),
.i_Sel(i_Sel[23])
);

Dummy_RO_cell D95(
.i_Enable(i_Enable),
.i_Sel(i_Sel[23])
);

Dummy_RO_cell D96(
.i_Enable(i_Enable),
.i_Sel(i_Sel[24])
);

Dummy_RO_cell D97(
.i_Enable(i_Enable),
.i_Sel(i_Sel[24])
);

Dummy_RO_cell D98(
.i_Enable(i_Enable),
.i_Sel(i_Sel[24])
);

Dummy_RO_cell D99(
.i_Enable(i_Enable),
.i_Sel(i_Sel[24])
);

Dummy_RO_cell D100(
.i_Enable(i_Enable),
.i_Sel(i_Sel[25])
);

Dummy_RO_cell D101(
.i_Enable(i_Enable),
.i_Sel(i_Sel[25])
);

Dummy_RO_cell D102(
.i_Enable(i_Enable),
.i_Sel(i_Sel[25])
);

Dummy_RO_cell D103(
.i_Enable(i_Enable),
.i_Sel(i_Sel[25])
);

Dummy_RO_cell D104(
.i_Enable(i_Enable),
.i_Sel(i_Sel[26])
);

Dummy_RO_cell D105(
.i_Enable(i_Enable),
.i_Sel(i_Sel[26])
);

Dummy_RO_cell D106(
.i_Enable(i_Enable),
.i_Sel(i_Sel[26])
);

Dummy_RO_cell D107(
.i_Enable(i_Enable),
.i_Sel(i_Sel[26])
);

Dummy_RO_cell D108(
.i_Enable(i_Enable),
.i_Sel(i_Sel[27])
);

Dummy_RO_cell D109(
.i_Enable(i_Enable),
.i_Sel(i_Sel[27])
);

Dummy_RO_cell D110(
.i_Enable(i_Enable),
.i_Sel(i_Sel[27])
);

Dummy_RO_cell D111(
.i_Enable(i_Enable),
.i_Sel(i_Sel[27])
);

Dummy_RO_cell D112(
.i_Enable(i_Enable),
.i_Sel(i_Sel[28])
);

Dummy_RO_cell D113(
.i_Enable(i_Enable),
.i_Sel(i_Sel[28])
);

Dummy_RO_cell D114(
.i_Enable(i_Enable),
.i_Sel(i_Sel[28])
);

Dummy_RO_cell D115(
.i_Enable(i_Enable),
.i_Sel(i_Sel[28])
);

Dummy_RO_cell D116(
.i_Enable(i_Enable),
.i_Sel(i_Sel[29])
);

Dummy_RO_cell D117(
.i_Enable(i_Enable),
.i_Sel(i_Sel[29])
);

Dummy_RO_cell D118(
.i_Enable(i_Enable),
.i_Sel(i_Sel[29])
);

Dummy_RO_cell D119(
.i_Enable(i_Enable),
.i_Sel(i_Sel[29])
);

Dummy_RO_cell D120(
.i_Enable(i_Enable),
.i_Sel(i_Sel[30])
);

Dummy_RO_cell D121(
.i_Enable(i_Enable),
.i_Sel(i_Sel[30])
);

Dummy_RO_cell D122(
.i_Enable(i_Enable),
.i_Sel(i_Sel[30])
);

Dummy_RO_cell D123(
.i_Enable(i_Enable),
.i_Sel(i_Sel[30])
);

Dummy_RO_cell D124(
.i_Enable(i_Enable),
.i_Sel(i_Sel[31])
);

Dummy_RO_cell D125(
.i_Enable(i_Enable),
.i_Sel(i_Sel[31])
);

Dummy_RO_cell D126(
.i_Enable(i_Enable),
.i_Sel(i_Sel[31])
);

Dummy_RO_cell D127(
.i_Enable(i_Enable),
.i_Sel(i_Sel[31])
);

endmodule 

